library verilog;
use verilog.vl_types.all;
entity DataMemory_vlg_vec_tst is
end DataMemory_vlg_vec_tst;
