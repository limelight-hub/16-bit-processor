library verilog;
use verilog.vl_types.all;
entity ram_vlg_vec_tst is
end ram_vlg_vec_tst;
