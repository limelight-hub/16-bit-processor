library verilog;
use verilog.vl_types.all;
entity ram4x4complete_vlg_vec_tst is
end ram4x4complete_vlg_vec_tst;
