library verilog;
use verilog.vl_types.all;
entity DMem64x16_vlg_vec_tst is
end DMem64x16_vlg_vec_tst;
