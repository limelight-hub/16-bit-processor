library verilog;
use verilog.vl_types.all;
entity stack4x4_vlg_vec_tst is
end stack4x4_vlg_vec_tst;
