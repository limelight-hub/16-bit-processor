library verilog;
use verilog.vl_types.all;
entity queue4x4_vlg_vec_tst is
end queue4x4_vlg_vec_tst;
