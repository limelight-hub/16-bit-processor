library verilog;
use verilog.vl_types.all;
entity ram_4x4_vlg_vec_tst is
end ram_4x4_vlg_vec_tst;
