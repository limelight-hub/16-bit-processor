library verilog;
use verilog.vl_types.all;
entity DMem_vlg_vec_tst is
end DMem_vlg_vec_tst;
